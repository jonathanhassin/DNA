
module deletion_restore #(
    parameter N = 100  // Number of digits in the word (will be set to 100)
)(
    input [2*N1-1:0] word_in,
    output logic [2*(N1+1)-1:0] word_out
);
    
	logic [] word_sum;
	logic [] diff_word;
	logic [] delta;
	logic [] gamma;
	
	
	
    diff_word diff_del_res (
	)
    
endmodule



